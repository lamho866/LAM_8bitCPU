module IM(
    input               clk,
    input               rst,
    input      [ 7:0]   PC_in,
    output     [15:0]   inst
);
parameter IM_DEPTH = 256;

reg [15:0] inst_mem[IM_DEPTH - 1:0];
assign inst = inst_mem[PC_in];
always @(posedge clk or posedge rst) begin
    if (rst) begin
        inst_mem[16'h0000] = 16'b001_11_010_000_00010;
        inst_mem[16'h0001] = 16'b001_11_011_000_00011;
        inst_mem[16'h0002] = 16'b001_11_100_000_00100;
        inst_mem[16'h0003] = 16'b001_11_111_000_00111;
        inst_mem[16'h0004] = 16'b000_00_010_010_011_00;
        inst_mem[16'h0005] = 16'b000_00_111_111_010_01;
        inst_mem[16'h0006] = 16'b000_00_011_011_100_10;
        inst_mem[16'h0007] = 16'b001_11_101_000_00101;
        inst_mem[16'h0008] = 16'b001_11_110_000_00110;
        inst_mem[16'h0009] = 16'b000_01_001_101_110_00;
        inst_mem[16'h000a] = 16'b000_01_001_010_111_01;
        inst_mem[16'h000b] = 16'b001_11_001_000_00001;
        inst_mem[16'h000c] = 16'b001_11_101_001_00100;
        inst_mem[16'h000d] = 16'b001_11_110_001_00011;
        inst_mem[16'h000e] = 16'b000_10_001_001_101_00;
        inst_mem[16'h000f] = 16'b000_10_001_001_110_01;
        inst_mem[16'h0010] = 16'b001_11_001_001_00011;
        inst_mem[16'h0011] = 16'b001_00_001_001_01100;
        inst_mem[16'h0012] = 16'b001_01_001_001_00011;
        inst_mem[16'h0013] = 16'b001_10_001_001_00011;
        inst_mem[16'h0014] = 16'b100_01_000000_001_00;
        inst_mem[16'h0015] = 16'b100_01_000000_010_01;
        inst_mem[16'h0016] = 16'b100_01_000000_011_10;
        inst_mem[16'h0017] = 16'b001_11_001_000_00000;
        inst_mem[16'h0018] = 16'b001_11_010_000_00000;
        inst_mem[16'h0019] = 16'b001_11_011_000_00000;
        inst_mem[16'h001a] = 16'b100_00_001_00000000;
        inst_mem[16'h001b] = 16'b100_00_010_00000001;
        inst_mem[16'h001c] = 16'b100_00_011_00000010;
        inst_mem[16'h001d] = 16'b000_00_000_000_001_00;
        inst_mem[16'h001e] = 16'b000_00_000_000_010_00;
        inst_mem[16'h001f] = 16'b000_00_000_000_011_00;
        inst_mem[16'h0020] = 16'b000_00_000_000_000_00;
    end else begin
        
    end
end
endmodule

